LIBRARY IEEE;
USE ieee.std_logic_1164.all;
--------------------------------------
ENTITY Bit8Mux16_1 IS

	PORT(	X1		:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X2		:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X3		:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X4		:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X5		:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X6		:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X7		:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X8		:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X9		:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X10	:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X11	:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X12	:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X13	:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X14	:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X15	:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			X16	:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
			sel	:	IN		STD_LOGIC_VECTOR(3 DOWNTO 0);
			Y		:	OUT	STD_LOGIC_VECTOR(7 DOWNTO 0));
			
END ENTITY Bit8Mux16_1;
--------------------------------------
ARCHITECTURE functional OF Bit8Mux16_1 IS
--------------------------------------
BEGIN

	WITH sel SELECT
		Y	<=	X1		WHEN	"0000",
				X2		WHEN	"0001",
				X3		WHEN	"0010",
				X4		WHEN	"0011",
				X5		WHEN	"0100",
				X6		WHEN	"0101",
				X7		WHEN	"0110",
				X8		WHEN	"0111",
				X9		WHEN	"1000",
				X10	WHEN	"1001",
				X11	WHEN	"1010",
				X12	WHEN	"1011",
				X13	WHEN	"1100",
				X14	WHEN	"1101",
				X15	WHEN	"1110",
				X16	WHEN	OTHERS;
	
END ARCHITECTURE	functional;